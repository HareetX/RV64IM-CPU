`include "defines.v"

module rom_top #(
    parameter BASE_IDX = `CPU_PC_RST_IDX,
    parameter IDX_LEN  = `CPU_PC_SIZE,
    parameter DATA_LEN = `CPU_INSTR_SIZE
) (
    input  [IDX_LEN-1:0]  rom_idx_i,
    output [DATA_LEN-1:0] rom_data_o,

    input  clk,
    input  rst_n
);

wire [IDX_LEN-1:0] rom_idx;

assign rom_idx = rom_idx_i - BASE_IDX;

rom_uninit #(`ROM_DATA_NUM, `ROM_DATA_IDXLEN, DATA_LEN) u_rom_uninit(
    .rom_idx_i   (rom_idx[`ROM_DATA_IDXLEN-1:0]   ),
    .rom_data_o  (rom_data_o                      ),
    .init_data_i ({
        32'h00000293,
        32'h00000313,
        32'hFFFFF3B7,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h16030A63,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h02038263,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h16039A63,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h18031263,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h1663CA63,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h18734263,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h16035A63,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h18735263,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h1803DA63,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h18736263,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h1863EA63,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h1863F263,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h18737A63,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000067,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE91FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hEA1FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE91FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hEA1FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE91FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hEA1FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE91FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE81FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE91FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE81FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE91FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00128293,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE81FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'hE91FF06F,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        32'h00000013,
        2048'd0
    } ), // 32-bit instructions
    .clk         (clk                              ),
    .rst_n       (rst_n                            )
);

endmodule