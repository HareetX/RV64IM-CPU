`include "defines.v"

module rom_top #(
    parameter BASE_IDX = `CPU_PC_RST_IDX,
    parameter IDX_LEN  = `CPU_PC_SIZE,
    parameter DATA_LEN = `CPU_INSTR_SIZE
) (
    input  [IDX_LEN-1:0]  rom_idx_i,
    output [DATA_LEN-1:0] rom_data_o,

    input  clk,
    input  rst_n
);

wire [IDX_LEN-1:0] rom_idx;

assign rom_idx = rom_idx_i - BASE_IDX;

rom_uninit #(`ROM_DATA_NUM, `ROM_DATA_IDXLEN, DATA_LEN) u_rom_uninit(
    .rom_idx_i   (rom_idx[`ROM_DATA_IDXLEN-1:0]   ),
    .rom_data_o  (rom_data_o                      ),
    .init_data_i ({
        32'b0000000_00001_00000_000_00001_0010011, // addi x1  x0  1 (00100093)
        32'b0000000_00001_00000_000_00010_0010011, // addi x2  x0  1 (00100113)
        32'b0000000_00001_00011_000_00000_0010011, // addi x0  x3  1
        32'b0000000_00010_00001_000_00011_0010011, // addi x3  x1  2
        32'b0000000_00010_00010_000_00100_0010011, // addi x4  x2  2
        32'b0000000_00010_00101_000_00000_0010011, // addi x0  x5  2

        32'b0100000_00011_00000_000_00101_0110011, // sub  x5  x0  x3
        32'b0000000_00100_00011_000_00110_0110011, // add  x6  x3  x4
        32'b0000000_00100_00011_000_00000_0110011, // add  x0  x3  x4

        32'b0000001_00011_00101_000_00111_0110011, // mul   x7  x5  x3
        32'b0000001_00110_00101_001_01000_0110011, // mulh  x8  x5  x6
        32'b0000001_00110_00101_010_01001_0110011, // mulsu x9  x5  x6
        32'b0000001_00101_00110_010_01010_0110011, // mulsu x10 x6  x5
        32'b0000001_00110_00101_011_01011_0110011, // mulu  x11 x5  x6

        32'b0000001_00011_00101_100_01100_0110011, // div   x12 x5  x3
        32'b0000001_00011_00101_101_01101_0110011, // divu  x13 x5  x3

        32'b0000001_00011_00101_110_01110_0110011, // rem   x14 x5  x3
        32'b0000001_00011_00101_111_01111_0110011, // remu  x15 x5  x3

        32'b0000000_00110_00011_011_10000_0110011, // sltu  x16 x3 x6
        32'b0000000_00000_00110_011_10001_0110011, // sltu  x17 x6 x0
        32'b0000000_00011_00011_011_10010_0110011, // sltu  x18 x3 x3

        32'b1111111_11111_00011_010_10011_0010011, // slti  x19 x3 -1
        32'b0000000_00110_00011_010_10100_0010011, // slti  x20 x3 6
        32'b0000000_00011_00011_010_10101_0010011, // slti  x21 x3 3

        32'b1111111_11111_00011_011_10110_0010011, // sltiu x22 x3 -1
        32'b0000000_00010_00011_011_10111_0010011, // sltiu x23 x3 2
        32'b0000000_00011_00011_011_11000_0010011, // sltiu x24 x3 3

        32'b0000000_00000_00000_000_00000_0000000,
        32'b0000000_00000_00000_000_00000_0000000,
        32'b0000000_00000_00000_000_00000_0000000,
        32'b0000000_00000_00000_000_00000_0000000,
        32'b0000000_00000_00000_000_00000_0000000
    } ), // 32-bit instructions
    .clk         (clk                              ),
    .rst_n       (rst_n                            )
);

endmodule