`include "defines.v"

module rom_top #(
    parameter BASE_IDX = `CPU_PC_RST_IDX,
    parameter IDX_LEN  = `CPU_PC_SIZE,
    parameter DATA_LEN = `CPU_INSTR_SIZE
) (
    input  [IDX_LEN-1:0]  rom_idx_i,
    output [DATA_LEN-1:0] rom_data_o,

    input  clk,
    input  rst_n
);

wire [IDX_LEN-1:0] rom_idx;

assign rom_idx = rom_idx_i - BASE_IDX;

rom_uninit #(`ROM_DATA_NUM, `ROM_DATA_IDXLEN, DATA_LEN) u_rom_uninit(
    .rom_idx_i   (rom_idx[`ROM_DATA_IDXLEN-1:0]   ),
    .rom_data_o  (rom_data_o                      ),
    .init_data_i ({
        32'b0000000_00001_00000_000_00001_0010011, // addi x1  x0  1
        32'b0000000_00001_00000_000_00010_0010011, // addi x2  x0  1
        32'b0000000_00001_00011_000_00000_0010011, // addi x0  x3  1
        32'b0000000_00010_00001_000_00011_0010011, // addi x3  x1  2
        32'b0000000_00010_00010_000_00100_0010011, // addi x4  x2  2
        32'b0000000_00010_00101_000_00000_0010011, // addi x0  x5  2
        32'b0000000_00011_00000_000_00101_0110011, // add  x5  x0  x
        32'b0000000_00100_00011_000_00110_0110011, // add  x6  x3  x
        32'b0000000_00100_00011_000_00000_0110011, // add  x0  x3  x
        32'b0100000_00000_00101_000_00111_0110011, // sub  x7  x5  x
        32'b0100000_00101_00110_000_01000_0110011, // sub  x8  x6  x
        32'b0100000_00110_00101_000_00000_0110011, // sub  x0  x5  x
        32'b0100000_00111_00000_000_01001_0110011, // sub  x9  x0  x
        32'b0000000_00001_11111_111_01010_0110111, // lui    x10 511
        32'b0000000_00001_11111_111_00000_0110111, // lui    x0  511
        32'b0000000_00001_11111_111_01011_0010111, // auipc x11 511
        32'b0000000_00001_11111_111_00000_0010111, // auipc x0  511
        32'b0000000_00110_00011_100_01100_0110011, // xor  x12 x3 x6
        32'b0000000_01110_00011_100_01101_0010011, // xori x13 x3 16
        32'b0000000_00110_00011_110_01110_0110011, // or   x14 x3 x6
        32'b0000000_01110_00011_110_01111_0010011, // ori  x15 x3 16
        32'b0000000_00110_00011_111_10000_0110011, // and  x16 x3 x6
        32'b0000000_01110_00011_111_10001_0010011, // andi x17 x3 16
        288'd0
    } ), // 32-bit instructions
    .clk         (clk                              ),
    .rst_n       (rst_n                            )
);

endmodule